module multi_packed_array;
  logic [2:0][3:0][3:0] arr;
  initial begin
    arr=$random;
    foreach(arr[i,j,k]) begin
      $display("arr[%0d][%0d][%0d]=%b",i,j,k,arr[i][j][k]);
    end
 end
endmodule

/* OUTPUT:
# run -all
# arr[2][3][3]=0
# arr[2][3][2]=0
# arr[2][3][1]=0
# arr[2][3][0]=0
# arr[2][2][3]=0
# arr[2][2][2]=0
# arr[2][2][1]=0
# arr[2][2][0]=0
# arr[2][1][3]=0
# arr[2][1][2]=0
# arr[2][1][1]=0
# arr[2][1][0]=0
# arr[2][0][3]=0
# arr[2][0][2]=0
# arr[2][0][1]=0
# arr[2][0][0]=0
# arr[1][3][3]=0
# arr[1][3][2]=0
# arr[1][3][1]=0
# arr[1][3][0]=1
# arr[1][2][3]=0
# arr[1][2][2]=0
# arr[1][2][1]=1
# arr[1][2][0]=0
# arr[1][1][3]=0
# arr[1][1][2]=0
# arr[1][1][1]=0
# arr[1][1][0]=1
# arr[1][0][3]=0
# arr[1][0][2]=1
# arr[1][0][1]=0
# arr[1][0][0]=1
# arr[0][3][3]=0
# arr[0][3][2]=0
# arr[0][3][1]=1
# arr[0][3][0]=1
# arr[0][2][3]=0
# arr[0][2][2]=1
# arr[0][2][1]=0
# arr[0][2][0]=1
# arr[0][1][3]=0
# arr[0][1][2]=0
# arr[0][1][1]=1
# arr[0][1][0]=0
# arr[0][0][3]=0
# arr[0][0][2]=1
# arr[0][0][1]=0
# arr[0][0][0]=0
*/
